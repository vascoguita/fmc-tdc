-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for TDC DMA Channel Control Registers
---------------------------------------------------------------------------------------
-- File           : tdc_dma_channel_regs.vhd
-- Author         : auto-generated by wbgen2 from wbgen/tdc_dma_channel_regs.wb
-- Created        : Wed Jul 18 23:25:00 2018
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE wbgen/tdc_dma_channel_regs.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wishbone_pkg.all;

use work.TDMA_wbgen2_pkg.all;


entity tdc_dma_channel_wb is
port (
  rst_n_i                                  : in     std_logic;
  clk_sys_i                                : in     std_logic;
  slave_i                                  : in     t_wishbone_slave_in;
  slave_o                                  : out    t_wishbone_slave_out;
  int_o                                    : out    std_logic;
  regs_i                                   : in     t_TDMA_in_registers;
  regs_o                                   : out    t_TDMA_out_registers
);
end tdc_dma_channel_wb;

architecture syn of tdc_dma_channel_wb is

signal tdma_csr_enable_int                      : std_logic      ;
signal tdma_csr_irq_timeout_int                 : std_logic_vector(9 downto 0);
signal tdma_csr_burst_size_int                  : std_logic_vector(9 downto 0);
signal tdma_csr_switch_buffers_dly0             : std_logic      ;
signal tdma_csr_switch_buffers_int              : std_logic      ;
signal ack_sreg                                 : std_logic_vector(9 downto 0);
signal rddata_reg                               : std_logic_vector(31 downto 0);
signal wrdata_reg                               : std_logic_vector(31 downto 0);
signal bwsel_reg                                : std_logic_vector(3 downto 0);
signal rwaddr_reg                               : std_logic_vector(2 downto 0);
signal ack_in_progress                          : std_logic      ;
signal wr_int                                   : std_logic      ;
signal rd_int                                   : std_logic      ;
signal allones                                  : std_logic_vector(31 downto 0);
signal allzeros                                 : std_logic_vector(31 downto 0);

begin
-- Some internal signals assignments
wrdata_reg <= slave_i.dat;
--
-- Main register bank access process.
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then
    ack_sreg <= "0000000000";
    ack_in_progress <= '0';
    rddata_reg <= "00000000000000000000000000000000";
    tdma_csr_enable_int <= '0';
    tdma_csr_irq_timeout_int <= "0000000000";
    tdma_csr_burst_size_int <= "0000000000";
    tdma_csr_switch_buffers_int <= '0';
    regs_o.tdma_csr_done_load_o <= '0';
    regs_o.tdma_csr_overflow_load_o <= '0';
    regs_o.tdma_cur_base_load_o <= '0';
    regs_o.tdma_cur_size_size_load_o <= '0';
    regs_o.tdma_cur_size_valid_load_o <= '0';
    regs_o.tdma_next_base_load_o <= '0';
    regs_o.tdma_next_size_size_load_o <= '0';
    regs_o.tdma_next_size_valid_load_o <= '0';
  elsif rising_edge(clk_sys_i) then
-- advance the ACK generator shift register
    ack_sreg(8 downto 0) <= ack_sreg(9 downto 1);
    ack_sreg(9) <= '0';
    if (ack_in_progress = '1') then
      if (ack_sreg(0) = '1') then
        tdma_csr_switch_buffers_int <= '0';
        regs_o.tdma_csr_done_load_o <= '0';
        regs_o.tdma_csr_overflow_load_o <= '0';
        regs_o.tdma_cur_base_load_o <= '0';
        regs_o.tdma_cur_size_size_load_o <= '0';
        regs_o.tdma_cur_size_valid_load_o <= '0';
        regs_o.tdma_next_base_load_o <= '0';
        regs_o.tdma_next_size_size_load_o <= '0';
        regs_o.tdma_next_size_valid_load_o <= '0';
        ack_in_progress <= '0';
      else
        regs_o.tdma_csr_done_load_o <= '0';
        regs_o.tdma_csr_overflow_load_o <= '0';
        regs_o.tdma_cur_base_load_o <= '0';
        regs_o.tdma_cur_size_size_load_o <= '0';
        regs_o.tdma_cur_size_valid_load_o <= '0';
        regs_o.tdma_next_base_load_o <= '0';
        regs_o.tdma_next_size_size_load_o <= '0';
        regs_o.tdma_next_size_valid_load_o <= '0';
      end if;
    else
      if ((slave_i.cyc = '1') and (slave_i.stb = '1')) then
        case rwaddr_reg(2 downto 0) is
        when "000" =>
          if (slave_i.we = '1') then
            tdma_csr_enable_int <= wrdata_reg(0);
            tdma_csr_irq_timeout_int <= wrdata_reg(10 downto 1);
            tdma_csr_burst_size_int <= wrdata_reg(20 downto 11);
            tdma_csr_switch_buffers_int <= wrdata_reg(21);
            regs_o.tdma_csr_done_load_o <= '1';
            regs_o.tdma_csr_overflow_load_o <= '1';
          end if;
          rddata_reg(0) <= tdma_csr_enable_int;
          rddata_reg(10 downto 1) <= tdma_csr_irq_timeout_int;
          rddata_reg(20 downto 11) <= tdma_csr_burst_size_int;
          rddata_reg(21) <= '0';
          rddata_reg(22) <= regs_i.tdma_csr_done_i;
          rddata_reg(23) <= regs_i.tdma_csr_overflow_i;
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(2) <= '1';
          ack_in_progress <= '1';
        when "001" =>
          if (slave_i.we = '1') then
            regs_o.tdma_cur_base_load_o <= '1';
          end if;
          rddata_reg(31 downto 0) <= regs_i.tdma_cur_base_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "010" =>
          if (slave_i.we = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tdma_cur_count_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "011" =>
          if (slave_i.we = '1') then
            regs_o.tdma_cur_size_size_load_o <= '1';
            regs_o.tdma_cur_size_valid_load_o <= '1';
          end if;
          rddata_reg(29 downto 0) <= regs_i.tdma_cur_size_size_i;
          rddata_reg(30) <= regs_i.tdma_cur_size_valid_i;
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "100" =>
          if (slave_i.we = '1') then
            regs_o.tdma_next_base_load_o <= '1';
          end if;
          rddata_reg(31 downto 0) <= regs_i.tdma_next_base_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "101" =>
          if (slave_i.we = '1') then
            regs_o.tdma_next_size_size_load_o <= '1';
            regs_o.tdma_next_size_valid_load_o <= '1';
          end if;
          rddata_reg(29 downto 0) <= regs_i.tdma_next_size_size_i;
          rddata_reg(30) <= regs_i.tdma_next_size_valid_i;
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when others =>
-- prevent the slave from hanging the bus on invalid address
          ack_in_progress <= '1';
          ack_sreg(0) <= '1';
        end case;
      end if;
    end if;
  end if;
end process;


-- Drive the data output bus
slave_o.dat <= rddata_reg;
-- Enable DMA
regs_o.tdma_csr_enable_o <= tdma_csr_enable_int;
-- IRQ Timeout (ms)
regs_o.tdma_csr_irq_timeout_o <= tdma_csr_irq_timeout_int;
-- Burst size (timestamps)
regs_o.tdma_csr_burst_size_o <= tdma_csr_burst_size_int;
-- Switch buffers
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then
    tdma_csr_switch_buffers_dly0 <= '0';
    regs_o.tdma_csr_switch_buffers_o <= '0';
  elsif rising_edge(clk_sys_i) then
    tdma_csr_switch_buffers_dly0 <= tdma_csr_switch_buffers_int;
    regs_o.tdma_csr_switch_buffers_o <= tdma_csr_switch_buffers_int and (not tdma_csr_switch_buffers_dly0);
  end if;
end process;


-- DMA complete
regs_o.tdma_csr_done_o <= wrdata_reg(22);
-- DMA overflow
regs_o.tdma_csr_overflow_o <= wrdata_reg(23);
-- Base address
regs_o.tdma_cur_base_o <= wrdata_reg(31 downto 0);
-- Number of data samples in the buffer
-- Size (in transfers)
regs_o.tdma_cur_size_size_o <= wrdata_reg(29 downto 0);
-- Valid flag
regs_o.tdma_cur_size_valid_o <= wrdata_reg(30);
-- Base address
regs_o.tdma_next_base_o <= wrdata_reg(31 downto 0);
-- Size (in transfers)
regs_o.tdma_next_size_size_o <= wrdata_reg(29 downto 0);
-- Valid flag
regs_o.tdma_next_size_valid_o <= wrdata_reg(30);
rwaddr_reg <= slave_i.adr(4 downto 2);
slave_o.stall <= (not ack_sreg(0)) and (slave_i.stb and slave_i.cyc);
slave_o.err <= '0';
slave_o.rty <= '0';
-- ACK signal generation. Just pass the LSB of ACK counter.
slave_o.ack <= ack_sreg(0);
end syn;
