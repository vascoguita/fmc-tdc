-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for TDC Direct Readout WB Slave
---------------------------------------------------------------------------------------
-- File           : ../fmc_tdc_direct_readout_slave_pkg.vhd
-- Author         : auto-generated by wbgen2 from fmc_tdc_direct_readout_slave.wb
-- Created        : Wed Mar 24 09:22:15 2021
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE fmc_tdc_direct_readout_slave.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wbgen2_pkg.all;

package dr_wbgen2_pkg is
  
  
  -- Input registers (user design -> WB slave)
  
  type t_dr_in_registers is record
    fifo_wr_req_i                            : std_logic;
    fifo_seconds_i                           : std_logic_vector(31 downto 0);
    fifo_cycles_i                            : std_logic_vector(31 downto 0);
    fifo_bins_i                              : std_logic_vector(17 downto 0);
    fifo_edge_i                              : std_logic;
    fifo_channel_i                           : std_logic_vector(3 downto 0);
    status_i                                 : std_logic;
    end record;
  
  constant c_dr_in_registers_init_value: t_dr_in_registers := (
    fifo_wr_req_i => '0',
    fifo_seconds_i => (others => '0'),
    fifo_cycles_i => (others => '0'),
    fifo_bins_i => (others => '0'),
    fifo_edge_i => '0',
    fifo_channel_i => (others => '0'),
    status_i => '0'
    );
    
    -- Output registers (WB slave -> user design)
    
    type t_dr_out_registers is record
      fifo_wr_full_o                           : std_logic;
      fifo_wr_empty_o                          : std_logic;
      fifo_wr_usedw_o                          : std_logic_vector(7 downto 0);
      chan_enable_o                            : std_logic_vector(4 downto 0);
      dead_time_o                              : std_logic_vector(23 downto 0);
      end record;
    
    constant c_dr_out_registers_init_value: t_dr_out_registers := (
      fifo_wr_full_o => '0',
      fifo_wr_empty_o => '0',
      fifo_wr_usedw_o => (others => '0'),
      chan_enable_o => (others => '0'),
      dead_time_o => (others => '0')
      );
    function "or" (left, right: t_dr_in_registers) return t_dr_in_registers;
    function f_x_to_zero (x:std_logic) return std_logic;
    function f_x_to_zero (x:std_logic_vector) return std_logic_vector;
end package;

package body dr_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
if x = '1' then
return '1';
else
return '0';
end if;
end function;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
variable tmp: std_logic_vector(x'length-1 downto 0);
begin
for i in 0 to x'length-1 loop
if(x(i) = '1') then
tmp(i):= '1';
else
tmp(i):= '0';
end if; 
end loop; 
return tmp;
end function;
function "or" (left, right: t_dr_in_registers) return t_dr_in_registers is
variable tmp: t_dr_in_registers;
begin
tmp.fifo_wr_req_i := f_x_to_zero(left.fifo_wr_req_i) or f_x_to_zero(right.fifo_wr_req_i);
tmp.fifo_seconds_i := f_x_to_zero(left.fifo_seconds_i) or f_x_to_zero(right.fifo_seconds_i);
tmp.fifo_cycles_i := f_x_to_zero(left.fifo_cycles_i) or f_x_to_zero(right.fifo_cycles_i);
tmp.fifo_bins_i := f_x_to_zero(left.fifo_bins_i) or f_x_to_zero(right.fifo_bins_i);
tmp.fifo_edge_i := f_x_to_zero(left.fifo_edge_i) or f_x_to_zero(right.fifo_edge_i);
tmp.fifo_channel_i := f_x_to_zero(left.fifo_channel_i) or f_x_to_zero(right.fifo_channel_i);
tmp.status_i := f_x_to_zero(left.status_i) or f_x_to_zero(right.status_i);
return tmp;
end function;
end package body;
