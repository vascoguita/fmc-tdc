-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for Timestamp FIFO
---------------------------------------------------------------------------------------
-- File           : timestamp_fifo_wbgen2_pkg.vhd
-- Author         : auto-generated by wbgen2 from wbgen/timestamp_fifo_wb.wb
-- Created        : Sun Sep  2 15:37:55 2018
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE wbgen/timestamp_fifo_wb.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wbgen2_pkg.all;
use work.wishbone_pkg.all;

package tsf_wbgen2_pkg is


  -- Input registers (user design -> WB slave)

  type t_tsf_in_registers is record
    fifo_wr_req_i                            : std_logic;
    fifo_ts0_i                               : std_logic_vector(31 downto 0);
    fifo_ts1_i                               : std_logic_vector(31 downto 0);
    fifo_ts2_i                               : std_logic_vector(31 downto 0);
    fifo_ts3_i                               : std_logic_vector(31 downto 0);
    delta1_i                                 : std_logic_vector(31 downto 0);
    delta2_i                                 : std_logic_vector(31 downto 0);
    delta3_i                                 : std_logic_vector(31 downto 0);
    csr_delta_ready_i                        : std_logic;
  end record;

  constant c_tsf_in_registers_init_value: t_tsf_in_registers := (
    fifo_wr_req_i => '0',
    fifo_ts0_i => (others => '0'),
    fifo_ts1_i => (others => '0'),
    fifo_ts2_i => (others => '0'),
    fifo_ts3_i => (others => '0'),
    delta1_i => (others => '0'),
    delta2_i => (others => '0'),
    delta3_i => (others => '0'),
    csr_delta_ready_i => '0'
  );

  -- Output registers (WB slave -> user design)

  type t_tsf_out_registers is record
    fifo_wr_full_o                           : std_logic;
    fifo_wr_empty_o                          : std_logic;
    fifo_wr_usedw_o                          : std_logic_vector(5 downto 0);
    offset1_o                                : std_logic_vector(31 downto 0);
    offset2_o                                : std_logic_vector(31 downto 0);
    offset3_o                                : std_logic_vector(31 downto 0);
    csr_delta_read_o                         : std_logic;
    csr_rst_seq_o                            : std_logic;
    csr_delta_ref_o                          : std_logic_vector(2 downto 0);
    csr_raw_mode_o                           : std_logic;
  end record;

  constant c_tsf_out_registers_init_value: t_tsf_out_registers := (
    fifo_wr_full_o => '0',
    fifo_wr_empty_o => '0',
    fifo_wr_usedw_o => (others => '0'),
    offset1_o => (others => '0'),
    offset2_o => (others => '0'),
    offset3_o => (others => '0'),
    csr_delta_read_o => '0',
    csr_rst_seq_o => '0',
    csr_delta_ref_o => (others => '0'),
    csr_raw_mode_o => '0'
  );

function "or" (left, right: t_tsf_in_registers) return t_tsf_in_registers;
function f_x_to_zero (x:std_logic) return std_logic;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector;

component timestamp_fifo_wb is
  port (
    rst_n_i                                  : in     std_logic;
    clk_sys_i                                : in     std_logic;
    slave_i                                  : in     t_wishbone_slave_in;
    slave_o                                  : out    t_wishbone_slave_out;
    int_o                                    : out    std_logic;
    regs_i                                   : in     t_tsf_in_registers;
    regs_o                                   : out    t_tsf_out_registers
  );
end component;

end package;

package body tsf_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
  if x = '1' then
    return '1';
  else
    return '0';
  end if;
end function;

function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
  variable tmp: std_logic_vector(x'length-1 downto 0);
begin
  for i in 0 to x'length-1 loop
    if(x(i) = 'X' or x(i) = 'U') then
      tmp(i):= '0';
    else
      tmp(i):=x(i);
    end if;
  end loop;
  return tmp;
end function;

function "or" (left, right: t_tsf_in_registers) return t_tsf_in_registers is
  variable tmp: t_tsf_in_registers;
begin
  tmp.fifo_wr_req_i := f_x_to_zero(left.fifo_wr_req_i) or f_x_to_zero(right.fifo_wr_req_i);
  tmp.fifo_ts0_i := f_x_to_zero(left.fifo_ts0_i) or f_x_to_zero(right.fifo_ts0_i);
  tmp.fifo_ts1_i := f_x_to_zero(left.fifo_ts1_i) or f_x_to_zero(right.fifo_ts1_i);
  tmp.fifo_ts2_i := f_x_to_zero(left.fifo_ts2_i) or f_x_to_zero(right.fifo_ts2_i);
  tmp.fifo_ts3_i := f_x_to_zero(left.fifo_ts3_i) or f_x_to_zero(right.fifo_ts3_i);
  tmp.delta1_i := f_x_to_zero(left.delta1_i) or f_x_to_zero(right.delta1_i);
  tmp.delta2_i := f_x_to_zero(left.delta2_i) or f_x_to_zero(right.delta2_i);
  tmp.delta3_i := f_x_to_zero(left.delta3_i) or f_x_to_zero(right.delta3_i);
  tmp.csr_delta_ready_i := f_x_to_zero(left.csr_delta_ready_i) or f_x_to_zero(right.csr_delta_ready_i);
  return tmp;
end function;

end package body;
