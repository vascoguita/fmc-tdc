`define ADDR_TDC_EIC_EIC_IDR           6'h20
`define TDC_EIC_EIC_IDR_TDC_FIFO1_OFFSET 0
`define TDC_EIC_EIC_IDR_TDC_FIFO1 32'h00000001
`define TDC_EIC_EIC_IDR_TDC_FIFO2_OFFSET 1
`define TDC_EIC_EIC_IDR_TDC_FIFO2 32'h00000002
`define TDC_EIC_EIC_IDR_TDC_FIFO3_OFFSET 2
`define TDC_EIC_EIC_IDR_TDC_FIFO3 32'h00000004
`define TDC_EIC_EIC_IDR_TDC_FIFO4_OFFSET 3
`define TDC_EIC_EIC_IDR_TDC_FIFO4 32'h00000008
`define TDC_EIC_EIC_IDR_TDC_FIFO5_OFFSET 4
`define TDC_EIC_EIC_IDR_TDC_FIFO5 32'h00000010
`define TDC_EIC_EIC_IDR_TDC_DMA1_OFFSET 5
`define TDC_EIC_EIC_IDR_TDC_DMA1 32'h00000020
`define TDC_EIC_EIC_IDR_TDC_DMA2_OFFSET 6
`define TDC_EIC_EIC_IDR_TDC_DMA2 32'h00000040
`define TDC_EIC_EIC_IDR_TDC_DMA3_OFFSET 7
`define TDC_EIC_EIC_IDR_TDC_DMA3 32'h00000080
`define TDC_EIC_EIC_IDR_TDC_DMA4_OFFSET 8
`define TDC_EIC_EIC_IDR_TDC_DMA4 32'h00000100
`define TDC_EIC_EIC_IDR_TDC_DMA5_OFFSET 9
`define TDC_EIC_EIC_IDR_TDC_DMA5 32'h00000200
`define ADDR_TDC_EIC_EIC_IER           6'h24
`define TDC_EIC_EIC_IER_TDC_FIFO1_OFFSET 0
`define TDC_EIC_EIC_IER_TDC_FIFO1 32'h00000001
`define TDC_EIC_EIC_IER_TDC_FIFO2_OFFSET 1
`define TDC_EIC_EIC_IER_TDC_FIFO2 32'h00000002
`define TDC_EIC_EIC_IER_TDC_FIFO3_OFFSET 2
`define TDC_EIC_EIC_IER_TDC_FIFO3 32'h00000004
`define TDC_EIC_EIC_IER_TDC_FIFO4_OFFSET 3
`define TDC_EIC_EIC_IER_TDC_FIFO4 32'h00000008
`define TDC_EIC_EIC_IER_TDC_FIFO5_OFFSET 4
`define TDC_EIC_EIC_IER_TDC_FIFO5 32'h00000010
`define TDC_EIC_EIC_IER_TDC_DMA1_OFFSET 5
`define TDC_EIC_EIC_IER_TDC_DMA1 32'h00000020
`define TDC_EIC_EIC_IER_TDC_DMA2_OFFSET 6
`define TDC_EIC_EIC_IER_TDC_DMA2 32'h00000040
`define TDC_EIC_EIC_IER_TDC_DMA3_OFFSET 7
`define TDC_EIC_EIC_IER_TDC_DMA3 32'h00000080
`define TDC_EIC_EIC_IER_TDC_DMA4_OFFSET 8
`define TDC_EIC_EIC_IER_TDC_DMA4 32'h00000100
`define TDC_EIC_EIC_IER_TDC_DMA5_OFFSET 9
`define TDC_EIC_EIC_IER_TDC_DMA5 32'h00000200
`define ADDR_TDC_EIC_EIC_IMR           6'h28
`define TDC_EIC_EIC_IMR_TDC_FIFO1_OFFSET 0
`define TDC_EIC_EIC_IMR_TDC_FIFO1 32'h00000001
`define TDC_EIC_EIC_IMR_TDC_FIFO2_OFFSET 1
`define TDC_EIC_EIC_IMR_TDC_FIFO2 32'h00000002
`define TDC_EIC_EIC_IMR_TDC_FIFO3_OFFSET 2
`define TDC_EIC_EIC_IMR_TDC_FIFO3 32'h00000004
`define TDC_EIC_EIC_IMR_TDC_FIFO4_OFFSET 3
`define TDC_EIC_EIC_IMR_TDC_FIFO4 32'h00000008
`define TDC_EIC_EIC_IMR_TDC_FIFO5_OFFSET 4
`define TDC_EIC_EIC_IMR_TDC_FIFO5 32'h00000010
`define TDC_EIC_EIC_IMR_TDC_DMA1_OFFSET 5
`define TDC_EIC_EIC_IMR_TDC_DMA1 32'h00000020
`define TDC_EIC_EIC_IMR_TDC_DMA2_OFFSET 6
`define TDC_EIC_EIC_IMR_TDC_DMA2 32'h00000040
`define TDC_EIC_EIC_IMR_TDC_DMA3_OFFSET 7
`define TDC_EIC_EIC_IMR_TDC_DMA3 32'h00000080
`define TDC_EIC_EIC_IMR_TDC_DMA4_OFFSET 8
`define TDC_EIC_EIC_IMR_TDC_DMA4 32'h00000100
`define TDC_EIC_EIC_IMR_TDC_DMA5_OFFSET 9
`define TDC_EIC_EIC_IMR_TDC_DMA5 32'h00000200
`define ADDR_TDC_EIC_EIC_ISR           6'h2c
`define TDC_EIC_EIC_ISR_TDC_FIFO1_OFFSET 0
`define TDC_EIC_EIC_ISR_TDC_FIFO1 32'h00000001
`define TDC_EIC_EIC_ISR_TDC_FIFO2_OFFSET 1
`define TDC_EIC_EIC_ISR_TDC_FIFO2 32'h00000002
`define TDC_EIC_EIC_ISR_TDC_FIFO3_OFFSET 2
`define TDC_EIC_EIC_ISR_TDC_FIFO3 32'h00000004
`define TDC_EIC_EIC_ISR_TDC_FIFO4_OFFSET 3
`define TDC_EIC_EIC_ISR_TDC_FIFO4 32'h00000008
`define TDC_EIC_EIC_ISR_TDC_FIFO5_OFFSET 4
`define TDC_EIC_EIC_ISR_TDC_FIFO5 32'h00000010
`define TDC_EIC_EIC_ISR_TDC_DMA1_OFFSET 5
`define TDC_EIC_EIC_ISR_TDC_DMA1 32'h00000020
`define TDC_EIC_EIC_ISR_TDC_DMA2_OFFSET 6
`define TDC_EIC_EIC_ISR_TDC_DMA2 32'h00000040
`define TDC_EIC_EIC_ISR_TDC_DMA3_OFFSET 7
`define TDC_EIC_EIC_ISR_TDC_DMA3 32'h00000080
`define TDC_EIC_EIC_ISR_TDC_DMA4_OFFSET 8
`define TDC_EIC_EIC_ISR_TDC_DMA4 32'h00000100
`define TDC_EIC_EIC_ISR_TDC_DMA5_OFFSET 9
`define TDC_EIC_EIC_ISR_TDC_DMA5 32'h00000200
