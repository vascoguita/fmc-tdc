// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CERN-OHL-W-2.0+

`define ADDR_TSF_DELTA1                6'h0
`define ADDR_TSF_DELTA2                6'h4
`define ADDR_TSF_DELTA3                6'h8
`define ADDR_TSF_OFFSET1               6'hc
`define ADDR_TSF_OFFSET2               6'h10
`define ADDR_TSF_OFFSET3               6'h14
`define ADDR_TSF_CSR                   6'h18
`define TSF_CSR_DELTA_READY_OFFSET 0
`define TSF_CSR_DELTA_READY 32'h00000001
`define TSF_CSR_DELTA_READ_OFFSET 1
`define TSF_CSR_DELTA_READ 32'h00000002
`define TSF_CSR_RST_SEQ_OFFSET 2
`define TSF_CSR_RST_SEQ 32'h00000004
`define TSF_CSR_DELTA_REF_OFFSET 3
`define TSF_CSR_DELTA_REF 32'h00000038
`define TSF_CSR_RAW_MODE_OFFSET 6
`define TSF_CSR_RAW_MODE 32'h00000040
`define ADDR_TSF_FIFO_R0               6'h1c
`define TSF_FIFO_R0_TS0_OFFSET 0
`define TSF_FIFO_R0_TS0 32'hffffffff
`define ADDR_TSF_FIFO_R1               6'h20
`define TSF_FIFO_R1_TS1_OFFSET 0
`define TSF_FIFO_R1_TS1 32'hffffffff
`define ADDR_TSF_FIFO_R2               6'h24
`define TSF_FIFO_R2_TS2_OFFSET 0
`define TSF_FIFO_R2_TS2 32'hffffffff
`define ADDR_TSF_FIFO_R3               6'h28
`define TSF_FIFO_R3_TS3_OFFSET 0
`define TSF_FIFO_R3_TS3 32'hffffffff
`define ADDR_TSF_FIFO_CSR              6'h2c
`define TSF_FIFO_CSR_FULL_OFFSET 16
`define TSF_FIFO_CSR_FULL 32'h00010000
`define TSF_FIFO_CSR_EMPTY_OFFSET 17
`define TSF_FIFO_CSR_EMPTY 32'h00020000
`define TSF_FIFO_CSR_CLEAR_BUS_OFFSET 18
`define TSF_FIFO_CSR_CLEAR_BUS 32'h00040000
`define TSF_FIFO_CSR_USEDW_OFFSET 0
`define TSF_FIFO_CSR_USEDW 32'h0000003f
