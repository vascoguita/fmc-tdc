// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CERN-OHL-W-2.0+

`define ADDR_TDC_BUF_CSR               5'h0
`define TDC_BUF_CSR_ENABLE_OFFSET 0
`define TDC_BUF_CSR_ENABLE 32'h00000001
`define TDC_BUF_CSR_IRQ_TIMEOUT_OFFSET 1
`define TDC_BUF_CSR_IRQ_TIMEOUT 32'h000007fe
`define TDC_BUF_CSR_BURST_SIZE_OFFSET 11
`define TDC_BUF_CSR_BURST_SIZE 32'h001ff800
`define TDC_BUF_CSR_SWITCH_BUFFERS_OFFSET 21
`define TDC_BUF_CSR_SWITCH_BUFFERS 32'h00200000
`define TDC_BUF_CSR_DONE_OFFSET 22
`define TDC_BUF_CSR_DONE 32'h00400000
`define TDC_BUF_CSR_OVERFLOW_OFFSET 23
`define TDC_BUF_CSR_OVERFLOW 32'h00800000
`define ADDR_TDC_BUF_CUR_BASE          5'h4
`define ADDR_TDC_BUF_CUR_COUNT         5'h8
`define ADDR_TDC_BUF_CUR_SIZE          5'hc
`define TDC_BUF_CUR_SIZE_SIZE_OFFSET 0
`define TDC_BUF_CUR_SIZE_SIZE 32'h3fffffff
`define TDC_BUF_CUR_SIZE_VALID_OFFSET 30
`define TDC_BUF_CUR_SIZE_VALID 32'h40000000
`define ADDR_TDC_BUF_NEXT_BASE         5'h10
`define ADDR_TDC_BUF_NEXT_SIZE         5'h14
`define TDC_BUF_NEXT_SIZE_SIZE_OFFSET 0
`define TDC_BUF_NEXT_SIZE_SIZE 32'h3fffffff
`define TDC_BUF_NEXT_SIZE_VALID_OFFSET 30
`define TDC_BUF_NEXT_SIZE_VALID 32'h40000000
