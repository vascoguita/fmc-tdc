// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CC0-1.0

`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG0 8'h0
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG1 8'h4
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG2 8'h8
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG3 8'hc
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG4 8'h10
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG5 8'h14
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG6 8'h18
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG7 8'h1c
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG11 8'h2c
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG12 8'h30
`define ADDR_TDC_CORE_CSR_ACAM_CFG_REG14 8'h38
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG0 8'h40
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG1 8'h44
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG2 8'h48
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG3 8'h4c
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG4 8'h50
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG5 8'h54
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG6 8'h58
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG7 8'h5c
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG8 8'h60
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG9 8'h64
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG10 8'h68
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG11 8'h6c
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG12 8'h70
`define ADDR_TDC_CORE_CSR_ACAM_RD_CFG_REG14 8'h78
`define ADDR_TDC_CORE_CSR_STARTING_UTC 8'h80
`define ADDR_TDC_CORE_CSR_ENABLE       8'h84
`define TDC_CORE_CSR_ENABLE_CH1_TERM_OFFSET 0
`define TDC_CORE_CSR_ENABLE_CH1_TERM 32'h00000001
`define TDC_CORE_CSR_ENABLE_CH2_TERM_OFFSET 1
`define TDC_CORE_CSR_ENABLE_CH2_TERM 32'h00000002
`define TDC_CORE_CSR_ENABLE_CH3_TERM_OFFSET 2
`define TDC_CORE_CSR_ENABLE_CH3_TERM 32'h00000004
`define TDC_CORE_CSR_ENABLE_CH4_TERM_OFFSET 3
`define TDC_CORE_CSR_ENABLE_CH4_TERM 32'h00000008
`define TDC_CORE_CSR_ENABLE_CH5_TERM_OFFSET 4
`define TDC_CORE_CSR_ENABLE_CH5_TERM 32'h00000010
`define TDC_CORE_CSR_ENABLE_ACAM_ACQ_OFFSET 7
`define TDC_CORE_CSR_ENABLE_ACAM_ACQ 32'h00000080
`define ADDR_TDC_CORE_CSR_C000FFEE_BREAK 8'h8c
`define ADDR_TDC_CORE_CSR_IRQ_TSTAMP_THRESH 8'h90
`define ADDR_TDC_CORE_CSR_IRQ_TIME_THRESH 8'h94
`define ADDR_TDC_CORE_CSR_DAC_WORD     8'h98
`define ADDR_TDC_CORE_CSR_UTC          8'ha0
`define ADDR_TDC_CORE_CSR_CORE_STATUS  8'hac
`define ADDR_TDC_CORE_CSR_WR_STAT      8'hb0
`define TDC_CORE_CSR_WR_STAT_WITH_WR_CORE_OFFSET 0
`define TDC_CORE_CSR_WR_STAT_WITH_WR_CORE 32'h00000001
`define TDC_CORE_CSR_WR_STAT_LINK_UP_OFFSET 1
`define TDC_CORE_CSR_WR_STAT_LINK_UP 32'h00000002
`define TDC_CORE_CSR_WR_STAT_AUX_CLK_LOCKED_OFFSET 2
`define TDC_CORE_CSR_WR_STAT_AUX_CLK_LOCKED 32'h00000004
`define TDC_CORE_CSR_WR_STAT_TIME_VALID_OFFSET 3
`define TDC_CORE_CSR_WR_STAT_TIME_VALID 32'h00000008
`define TDC_CORE_CSR_WR_STAT_AUX_CLK_LOCK_EN_OFFSET 4
`define TDC_CORE_CSR_WR_STAT_AUX_CLK_LOCK_EN 32'h00000010
`define ADDR_TDC_CORE_CSR_WR_CTRL      8'hb4
`define TDC_CORE_CSR_WR_CTRL_EN_OFFSET 0
`define TDC_CORE_CSR_WR_CTRL_EN 32'h00000001
`define TDC_CORE_CSR_WR_CTRL_UNUSED_OFFSET 1
`define TDC_CORE_CSR_WR_CTRL_UNUSED 32'hfffffffe
`define ADDR_TDC_CORE_CSR_TEST0        8'hb8
`define TDC_CORE_CSR_TEST0_FAKE_TS_PERIOD_OFFSET 0
`define TDC_CORE_CSR_TEST0_FAKE_TS_PERIOD 32'h0fffffff
`define TDC_CORE_CSR_TEST0_FAKE_TS_CH_OFFSET 28
`define TDC_CORE_CSR_TEST0_FAKE_TS_CH 32'h70000000
`define TDC_CORE_CSR_TEST0_FAKE_TS_EN_OFFSET 31
`define TDC_CORE_CSR_TEST0_FAKE_TS_EN 32'h80000000
`define ADDR_TDC_CORE_CSR_TEST1        8'hbc
`define ADDR_TDC_CORE_CSR_CTRL         8'hfc
`define TDC_CORE_CSR_CTRL_ACTIVATE_ACQ_P_OFFSET 0
`define TDC_CORE_CSR_CTRL_ACTIVATE_ACQ_P 32'h00000001
`define TDC_CORE_CSR_CTRL_DEACTIVATE_ACQ_P_OFFSET 1
`define TDC_CORE_CSR_CTRL_DEACTIVATE_ACQ_P 32'h00000002
`define TDC_CORE_CSR_CTRL_LOAD_ACAM_CFG_P_OFFSET 2
`define TDC_CORE_CSR_CTRL_LOAD_ACAM_CFG_P 32'h00000004
`define TDC_CORE_CSR_CTRL_RD_ACAM_CFG_P_OFFSET 3
`define TDC_CORE_CSR_CTRL_RD_ACAM_CFG_P 32'h00000008
`define TDC_CORE_CSR_CTRL_RD_ACAM_STATUS_P_OFFSET 4
`define TDC_CORE_CSR_CTRL_RD_ACAM_STATUS_P 32'h00000010
`define TDC_CORE_CSR_CTRL_RD_ACAM_IFIFO1_P_OFFSET 5
`define TDC_CORE_CSR_CTRL_RD_ACAM_IFIFO1_P 32'h00000020
`define TDC_CORE_CSR_CTRL_RD_ACAM_IFIFO2_P_OFFSET 6
`define TDC_CORE_CSR_CTRL_RD_ACAM_IFIFO2_P 32'h00000040
`define TDC_CORE_CSR_CTRL_RD_ACAM_START01_P_OFFSET 7
`define TDC_CORE_CSR_CTRL_RD_ACAM_START01_P 32'h00000080
`define TDC_CORE_CSR_CTRL_RST_ACAM_P_OFFSET 8
`define TDC_CORE_CSR_CTRL_RST_ACAM_P 32'h00000100
`define TDC_CORE_CSR_CTRL_LOAD_UTC_P_OFFSET 9
`define TDC_CORE_CSR_CTRL_LOAD_UTC_P 32'h00000200
`define TDC_CORE_CSR_CTRL_LOAD_DAC_P_OFFSET 10
`define TDC_CORE_CSR_CTRL_LOAD_DAC_P 32'h00000400
