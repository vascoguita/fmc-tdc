// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CERN-OHL-W-2.0+

`define ADDR_DMA_CTRL                  6'h0
`define ADDR_DMA_STAT                  6'h4
`define ADDR_DMA_CSTART                6'h8
`define ADDR_DMA_HSTARTL               6'hc
`define ADDR_DMA_HSTARTH               6'h10
`define ADDR_DMA_LEN                   6'h14
`define ADDR_DMA_NEXTL                 6'h18
`define ADDR_DMA_NEXTH                 6'h1c
`define ADDR_DMA_ATTRIB                6'h20
