// SPDX-FileCopyrightText: 2022 CERN (home.cern)
//
// SPDX-License-Identifier: CC0-1.0

`define SPEC_BASE_REGS_SIZE 8192
`define ADDR_SPEC_BASE_REGS_METADATA 'h0
`define SPEC_BASE_REGS_METADATA_SIZE 64
`define ADDR_SPEC_BASE_REGS_CSR 'h40
`define SPEC_BASE_REGS_CSR_SIZE 32
`define ADDR_SPEC_BASE_REGS_CSR_APP_OFFSET 'h40
`define ADDR_SPEC_BASE_REGS_CSR_RESETS 'h44
`define SPEC_BASE_REGS_CSR_RESETS_GLOBAL_OFFSET 0
`define SPEC_BASE_REGS_CSR_RESETS_GLOBAL 'h1
`define SPEC_BASE_REGS_CSR_RESETS_APPL_OFFSET 1
`define SPEC_BASE_REGS_CSR_RESETS_APPL 'h2
`define ADDR_SPEC_BASE_REGS_CSR_FMC_PRESENCE 'h48
`define ADDR_SPEC_BASE_REGS_CSR_GN4124_STATUS 'h4c
`define ADDR_SPEC_BASE_REGS_CSR_DDR_STATUS 'h50
`define SPEC_BASE_REGS_CSR_DDR_STATUS_CALIB_DONE_OFFSET 0
`define SPEC_BASE_REGS_CSR_DDR_STATUS_CALIB_DONE 'h1
`define ADDR_SPEC_BASE_REGS_CSR_PCB_REV 'h54
`define SPEC_BASE_REGS_CSR_PCB_REV_REV_OFFSET 0
`define SPEC_BASE_REGS_CSR_PCB_REV_REV 'hf
`define ADDR_SPEC_BASE_REGS_THERM_ID 'h70
`define SPEC_BASE_REGS_THERM_ID_SIZE 16
`define ADDR_SPEC_BASE_REGS_FMC_I2C 'h80
`define SPEC_BASE_REGS_FMC_I2C_SIZE 32
`define ADDR_SPEC_BASE_REGS_FLASH_SPI 'ha0
`define SPEC_BASE_REGS_FLASH_SPI_SIZE 32
`define ADDR_SPEC_BASE_REGS_DMA 'hc0
`define SPEC_BASE_REGS_DMA_SIZE 64
`define ADDR_SPEC_BASE_REGS_VIC 'h100
`define SPEC_BASE_REGS_VIC_SIZE 256
`define ADDR_SPEC_BASE_REGS_BUILDINFO 'h200
`define SPEC_BASE_REGS_BUILDINFO_SIZE 256
`define ADDR_SPEC_BASE_REGS_WRC_REGS 'h1000
`define SPEC_BASE_REGS_WRC_REGS_SIZE 4096
