-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for TDC Onewire Master
---------------------------------------------------------------------------------------
-- File           : tdc_onewire_wb.vhd
-- Author         : auto-generated by wbgen2 from wbgen/tdc_onewire_wb.wb
-- Created        : Tue Sep 11 11:16:49 2018
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE wbgen/tdc_onewire_wb.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wishbone_pkg.all;

use work.TDC_OW_wbgen2_pkg.all;


entity tdc_onewire_wb is
port (
  rst_n_i                                  : in     std_logic;
  clk_sys_i                                : in     std_logic;
  slave_i                                  : in     t_wishbone_slave_in;
  slave_o                                  : out    t_wishbone_slave_out;
  int_o                                    : out    std_logic;
  regs_i                                   : in     t_TDC_OW_in_registers;
  regs_o                                   : out    t_TDC_OW_out_registers
);
end tdc_onewire_wb;

architecture syn of tdc_onewire_wb is

signal ack_sreg                                 : std_logic_vector(9 downto 0);
signal rddata_reg                               : std_logic_vector(31 downto 0);
signal wrdata_reg                               : std_logic_vector(31 downto 0);
signal bwsel_reg                                : std_logic_vector(3 downto 0);
signal rwaddr_reg                               : std_logic_vector(1 downto 0);
signal ack_in_progress                          : std_logic      ;
signal wr_int                                   : std_logic      ;
signal rd_int                                   : std_logic      ;
signal allones                                  : std_logic_vector(31 downto 0);
signal allzeros                                 : std_logic_vector(31 downto 0);

begin
-- Some internal signals assignments
wrdata_reg <= slave_i.dat;
-- 
-- Main register bank access process.
process (clk_sys_i, rst_n_i)
begin
  if (rst_n_i = '0') then 
    ack_sreg <= "0000000000";
    ack_in_progress <= '0';
    rddata_reg <= "00000000000000000000000000000000";
    regs_o.tdc_ow_csr_valid_load_o <= '0';
  elsif rising_edge(clk_sys_i) then
-- advance the ACK generator shift register
    ack_sreg(8 downto 0) <= ack_sreg(9 downto 1);
    ack_sreg(9) <= '0';
    if (ack_in_progress = '1') then
      if (ack_sreg(0) = '1') then
        regs_o.tdc_ow_csr_valid_load_o <= '0';
        ack_in_progress <= '0';
      else
        regs_o.tdc_ow_csr_valid_load_o <= '0';
      end if;
    else
      if ((slave_i.cyc = '1') and (slave_i.stb = '1')) then
        case rwaddr_reg(1 downto 0) is
        when "00" => 
          if (slave_i.we = '1') then
            regs_o.tdc_ow_csr_valid_load_o <= '1';
          end if;
          rddata_reg(0) <= regs_i.tdc_ow_csr_valid_i;
          rddata_reg(1) <= 'X';
          rddata_reg(2) <= 'X';
          rddata_reg(3) <= 'X';
          rddata_reg(4) <= 'X';
          rddata_reg(5) <= 'X';
          rddata_reg(6) <= 'X';
          rddata_reg(7) <= 'X';
          rddata_reg(8) <= 'X';
          rddata_reg(9) <= 'X';
          rddata_reg(10) <= 'X';
          rddata_reg(11) <= 'X';
          rddata_reg(12) <= 'X';
          rddata_reg(13) <= 'X';
          rddata_reg(14) <= 'X';
          rddata_reg(15) <= 'X';
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "01" => 
          if (slave_i.we = '1') then
          end if;
          rddata_reg(15 downto 0) <= regs_i.tdc_ow_temp_i;
          rddata_reg(16) <= 'X';
          rddata_reg(17) <= 'X';
          rddata_reg(18) <= 'X';
          rddata_reg(19) <= 'X';
          rddata_reg(20) <= 'X';
          rddata_reg(21) <= 'X';
          rddata_reg(22) <= 'X';
          rddata_reg(23) <= 'X';
          rddata_reg(24) <= 'X';
          rddata_reg(25) <= 'X';
          rddata_reg(26) <= 'X';
          rddata_reg(27) <= 'X';
          rddata_reg(28) <= 'X';
          rddata_reg(29) <= 'X';
          rddata_reg(30) <= 'X';
          rddata_reg(31) <= 'X';
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "10" => 
          if (slave_i.we = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tdc_ow_id_h_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when "11" => 
          if (slave_i.we = '1') then
          end if;
          rddata_reg(31 downto 0) <= regs_i.tdc_ow_id_l_i;
          ack_sreg(0) <= '1';
          ack_in_progress <= '1';
        when others =>
-- prevent the slave from hanging the bus on invalid address
          ack_in_progress <= '1';
          ack_sreg(0) <= '1';
        end case;
      end if;
    end if;
  end if;
end process;


-- Drive the data output bus
slave_o.dat <= rddata_reg;
-- Temperature & ID valid
regs_o.tdc_ow_csr_valid_o <= wrdata_reg(0);
-- Temperature
-- Unique ID (32 highest bits)
-- Unique ID (32 lowest bits)
rwaddr_reg <= slave_i.adr(3 downto 2);
slave_o.stall <= (not ack_sreg(0)) and (slave_i.stb and slave_i.cyc);
slave_o.err <= '0';
slave_o.rty <= '0';
-- ACK signal generation. Just pass the LSB of ACK counter.
slave_o.ack <= ack_sreg(0);
end syn;
