-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for TDC DMA Channel Control Registers
---------------------------------------------------------------------------------------
-- File           : tdc_dma_channel_wbgen2_pkg.vhd
-- Author         : auto-generated by wbgen2 from wbgen/tdc_dma_channel_regs.wb
-- Created        : Wed Jul 18 23:25:00 2018
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE wbgen/tdc_dma_channel_regs.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wishbone_pkg.all;

package TDMA_wbgen2_pkg is


  -- Input registers (user design -> WB slave)

  type t_TDMA_in_registers is record
    tdma_csr_done_i                          : std_logic;
    tdma_csr_overflow_i                      : std_logic;
    tdma_cur_base_i                          : std_logic_vector(31 downto 0);
    tdma_cur_count_i                         : std_logic_vector(31 downto 0);
    tdma_cur_size_size_i                     : std_logic_vector(29 downto 0);
    tdma_cur_size_valid_i                    : std_logic;
    tdma_next_base_i                         : std_logic_vector(31 downto 0);
    tdma_next_size_size_i                    : std_logic_vector(29 downto 0);
    tdma_next_size_valid_i                   : std_logic;
  end record;

  constant c_TDMA_in_registers_init_value: t_TDMA_in_registers := (
    tdma_csr_done_i => '0',
    tdma_csr_overflow_i => '0',
    tdma_cur_base_i => (others => '0'),
    tdma_cur_count_i => (others => '0'),
    tdma_cur_size_size_i => (others => '0'),
    tdma_cur_size_valid_i => '0',
    tdma_next_base_i => (others => '0'),
    tdma_next_size_size_i => (others => '0'),
    tdma_next_size_valid_i => '0'
  );

  -- Output registers (WB slave -> user design)

  type t_TDMA_out_registers is record
    tdma_csr_enable_o                        : std_logic;
    tdma_csr_irq_timeout_o                   : std_logic_vector(9 downto 0);
    tdma_csr_burst_size_o                    : std_logic_vector(9 downto 0);
    tdma_csr_switch_buffers_o                : std_logic;
    tdma_csr_done_o                          : std_logic;
    tdma_csr_done_load_o                     : std_logic;
    tdma_csr_overflow_o                      : std_logic;
    tdma_csr_overflow_load_o                 : std_logic;
    tdma_cur_base_o                          : std_logic_vector(31 downto 0);
    tdma_cur_base_load_o                     : std_logic;
    tdma_cur_size_size_o                     : std_logic_vector(29 downto 0);
    tdma_cur_size_size_load_o                : std_logic;
    tdma_cur_size_valid_o                    : std_logic;
    tdma_cur_size_valid_load_o               : std_logic;
    tdma_next_base_o                         : std_logic_vector(31 downto 0);
    tdma_next_base_load_o                    : std_logic;
    tdma_next_size_size_o                    : std_logic_vector(29 downto 0);
    tdma_next_size_size_load_o               : std_logic;
    tdma_next_size_valid_o                   : std_logic;
    tdma_next_size_valid_load_o              : std_logic;
  end record;

  constant c_TDMA_out_registers_init_value: t_TDMA_out_registers := (
    tdma_csr_enable_o => '0',
    tdma_csr_irq_timeout_o => (others => '0'),
    tdma_csr_burst_size_o => (others => '0'),
    tdma_csr_switch_buffers_o => '0',
    tdma_csr_done_o => '0',
    tdma_csr_done_load_o => '0',
    tdma_csr_overflow_o => '0',
    tdma_csr_overflow_load_o => '0',
    tdma_cur_base_o => (others => '0'),
    tdma_cur_base_load_o => '0',
    tdma_cur_size_size_o => (others => '0'),
    tdma_cur_size_size_load_o => '0',
    tdma_cur_size_valid_o => '0',
    tdma_cur_size_valid_load_o => '0',
    tdma_next_base_o => (others => '0'),
    tdma_next_base_load_o => '0',
    tdma_next_size_size_o => (others => '0'),
    tdma_next_size_size_load_o => '0',
    tdma_next_size_valid_o => '0',
    tdma_next_size_valid_load_o => '0'
  );

function "or" (left, right: t_TDMA_in_registers) return t_TDMA_in_registers;
function f_x_to_zero (x:std_logic) return std_logic;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector;

component tdc_dma_channel_wb is
  port (
    rst_n_i                                  : in     std_logic;
    clk_sys_i                                : in     std_logic;
    slave_i                                  : in     t_wishbone_slave_in;
    slave_o                                  : out    t_wishbone_slave_out;
    int_o                                    : out    std_logic;
    regs_i                                   : in     t_TDMA_in_registers;
    regs_o                                   : out    t_TDMA_out_registers
  );
end component;

end package;

package body TDMA_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
  if x = '1' then
    return '1';
  else
    return '0';
  end if;
end function;

function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
  variable tmp: std_logic_vector(x'length-1 downto 0);
begin
  for i in 0 to x'length-1 loop
    if(x(i) = 'X' or x(i) = 'U') then
      tmp(i):= '0';
    else
      tmp(i):=x(i);
    end if;
  end loop;
  return tmp;
end function;

function "or" (left, right: t_TDMA_in_registers) return t_TDMA_in_registers is
  variable tmp: t_TDMA_in_registers;
begin
  tmp.tdma_csr_done_i := f_x_to_zero(left.tdma_csr_done_i) or f_x_to_zero(right.tdma_csr_done_i);
  tmp.tdma_csr_overflow_i := f_x_to_zero(left.tdma_csr_overflow_i) or f_x_to_zero(right.tdma_csr_overflow_i);
  tmp.tdma_cur_base_i := f_x_to_zero(left.tdma_cur_base_i) or f_x_to_zero(right.tdma_cur_base_i);
  tmp.tdma_cur_count_i := f_x_to_zero(left.tdma_cur_count_i) or f_x_to_zero(right.tdma_cur_count_i);
  tmp.tdma_cur_size_size_i := f_x_to_zero(left.tdma_cur_size_size_i) or f_x_to_zero(right.tdma_cur_size_size_i);
  tmp.tdma_cur_size_valid_i := f_x_to_zero(left.tdma_cur_size_valid_i) or f_x_to_zero(right.tdma_cur_size_valid_i);
  tmp.tdma_next_base_i := f_x_to_zero(left.tdma_next_base_i) or f_x_to_zero(right.tdma_next_base_i);
  tmp.tdma_next_size_size_i := f_x_to_zero(left.tdma_next_size_size_i) or f_x_to_zero(right.tdma_next_size_size_i);
  tmp.tdma_next_size_valid_i := f_x_to_zero(left.tdma_next_size_valid_i) or f_x_to_zero(right.tdma_next_size_valid_i);
  return tmp;
end function;

end package body;
