-- SPDX-FileCopyrightText: 2022 CERN (home.cern)
--
-- SPDX-License-Identifier: CERN-OHL-W-2.0+

---------------------------------------------------------------------------------------
-- Title          : Wishbone slave core for TDC Onewire Master
---------------------------------------------------------------------------------------
-- File           : tdc_onewire_wbgen2_pkg.vhd
-- Author         : auto-generated by wbgen2 from wbgen/tdc_onewire_wb.wb
-- Created        : Tue Sep 11 11:16:49 2018
-- Standard       : VHDL'87
---------------------------------------------------------------------------------------
-- THIS FILE WAS GENERATED BY wbgen2 FROM SOURCE FILE wbgen/tdc_onewire_wb.wb
-- DO NOT HAND-EDIT UNLESS IT'S ABSOLUTELY NECESSARY!
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.wishbone_pkg.all;

package TDC_OW_wbgen2_pkg is
  
  
  -- Input registers (user design -> WB slave)
  
  type t_TDC_OW_in_registers is record
    tdc_ow_csr_valid_i                       : std_logic;
    tdc_ow_temp_i                            : std_logic_vector(15 downto 0);
    tdc_ow_id_h_i                            : std_logic_vector(31 downto 0);
    tdc_ow_id_l_i                            : std_logic_vector(31 downto 0);
  end record;
  
  constant c_TDC_OW_in_registers_init_value: t_TDC_OW_in_registers := (
    tdc_ow_csr_valid_i => '0',
    tdc_ow_temp_i => (others => '0'),
    tdc_ow_id_h_i => (others => '0'),
    tdc_ow_id_l_i => (others => '0')
  );
  
  -- Output registers (WB slave -> user design)
  
  type t_TDC_OW_out_registers is record
    tdc_ow_csr_valid_o                       : std_logic;
    tdc_ow_csr_valid_load_o                  : std_logic;
  end record;
  
  constant c_TDC_OW_out_registers_init_value: t_TDC_OW_out_registers := (
    tdc_ow_csr_valid_o => '0',
    tdc_ow_csr_valid_load_o => '0'
  );

function "or" (left, right: t_TDC_OW_in_registers) return t_TDC_OW_in_registers;
function f_x_to_zero (x:std_logic) return std_logic;
function f_x_to_zero (x:std_logic_vector) return std_logic_vector;

component tdc_onewire_wb is
  port (
    rst_n_i                                  : in     std_logic;
    clk_sys_i                                : in     std_logic;
    slave_i                                  : in     t_wishbone_slave_in;
    slave_o                                  : out    t_wishbone_slave_out;
    int_o                                    : out    std_logic;
    regs_i                                   : in     t_TDC_OW_in_registers;
    regs_o                                   : out    t_TDC_OW_out_registers
  );
end component;

end package;

package body TDC_OW_wbgen2_pkg is
function f_x_to_zero (x:std_logic) return std_logic is
begin
  if x = '1' then
    return '1';
  else
    return '0';
  end if;
end function;

function f_x_to_zero (x:std_logic_vector) return std_logic_vector is
  variable tmp: std_logic_vector(x'length-1 downto 0);
begin
  for i in 0 to x'length-1 loop
    if(x(i) = 'X' or x(i) = 'U') then
      tmp(i):= '0';
    else
      tmp(i):=x(i);
    end if; 
  end loop; 
  return tmp;
end function;

function "or" (left, right: t_TDC_OW_in_registers) return t_TDC_OW_in_registers is
  variable tmp: t_TDC_OW_in_registers;
begin
  tmp.tdc_ow_csr_valid_i := f_x_to_zero(left.tdc_ow_csr_valid_i) or f_x_to_zero(right.tdc_ow_csr_valid_i);
  tmp.tdc_ow_temp_i := f_x_to_zero(left.tdc_ow_temp_i) or f_x_to_zero(right.tdc_ow_temp_i);
  tmp.tdc_ow_id_h_i := f_x_to_zero(left.tdc_ow_id_h_i) or f_x_to_zero(right.tdc_ow_id_h_i);
  tmp.tdc_ow_id_l_i := f_x_to_zero(left.tdc_ow_id_l_i) or f_x_to_zero(right.tdc_ow_id_l_i);
  return tmp;
end function;

end package body;
